// hw_qsys.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module hw_qsys (
		input  wire        clk_clk,             //   clk.clk
		output wire        hdmi_clk_mm,         //  hdmi.clk_mm
		output wire        hdmi_clk_pix_p,      //      .clk_pix_p
		output wire        hdmi_clk_pix_n,      //      .clk_pix_n
		output wire        hdmi_red_p,          //      .red_p
		output wire        hdmi_red_n,          //      .red_n
		output wire        hdmi_green_p,        //      .green_p
		output wire        hdmi_green_n,        //      .green_n
		output wire        hdmi_blue_p,         //      .blue_p
		output wire        hdmi_blue_n,         //      .blue_n
		output wire [10:0] hdmi_x,              //      .x
		output wire [10:0] hdmi_y,              //      .y
		output wire [10:0] hdmi_horz,           //      .horz
		output wire [10:0] hdmi_vert,           //      .vert
		input  wire        reset_reset_n,       // reset.reset_n
		input  wire        slave_read,          // slave.read
		input  wire        slave_write,         //      .write
		input  wire [9:0]  slave_address,       //      .address
		input  wire [31:0] slave_writedata,     //      .writedata
		input  wire        slave_burstcount,    //      .burstcount
		input  wire [3:0]  slave_byteenable,    //      .byteenable
		output wire        slave_waitrequest,   //      .waitrequest
		output wire        slave_readdatavalid, //      .readdatavalid
		output wire [31:0] slave_readdata       //      .readdata
	);

	wire    altpll_0_c0_clk;                // altpll_0:c0 -> hdmi_mm_0:clk_x10
	wire    altpll_0_c1_clk;                // altpll_0:c1 -> [hdmi_mm_0:clk, rst_controller:clk]
	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> hdmi_mm_0:reset

	hw_qsys_altpll_0 altpll_0 (
		.clk                (clk_clk),         //       inclk_interface.clk
		.reset              (~reset_reset_n),  // inclk_interface_reset.reset
		.read               (),                //             pll_slave.read
		.write              (),                //                      .write
		.address            (),                //                      .address
		.readdata           (),                //                      .readdata
		.writedata          (),                //                      .writedata
		.c0                 (altpll_0_c0_clk), //                    c0.clk
		.c1                 (altpll_0_c1_clk), //                    c1.clk
		.scandone           (),                //           (terminated)
		.scandataout        (),                //           (terminated)
		.c2                 (),                //           (terminated)
		.c3                 (),                //           (terminated)
		.c4                 (),                //           (terminated)
		.areset             (1'b0),            //           (terminated)
		.locked             (),                //           (terminated)
		.phasedone          (),                //           (terminated)
		.phasecounterselect (3'b000),          //           (terminated)
		.phaseupdown        (1'b0),            //           (terminated)
		.phasestep          (1'b0),            //           (terminated)
		.scanclk            (1'b0),            //           (terminated)
		.scanclkena         (1'b0),            //           (terminated)
		.scandata           (1'b0),            //           (terminated)
		.configupdate       (1'b0)             //           (terminated)
	);

	hdmi_mm #(
		.horz_front_porch (18),
		.horz_sync        (60),
		.horz_back_porch  (112),
		.horz_pix         (1024),
		.vert_front_porch (18),
		.vert_sync        (60),
		.vert_back_porch  (112),
		.vert_pix         (600)
	) hdmi_mm_0 (
		.clk             (altpll_0_c1_clk),                //        clock.clk
		.reset           (rst_controller_reset_out_reset), //        reset.reset
		.clk_mm          (hdmi_clk_mm),                    //      hdmi_mm.clk_mm
		.clk_pix_p       (hdmi_clk_pix_p),                 //             .clk_pix_p
		.clk_pix_n       (hdmi_clk_pix_n),                 //             .clk_pix_n
		.red_p           (hdmi_red_p),                     //             .red_p
		.red_n           (hdmi_red_n),                     //             .red_n
		.green_p         (hdmi_green_p),                   //             .green_p
		.green_n         (hdmi_green_n),                   //             .green_n
		.blue_p          (hdmi_blue_p),                    //             .blue_p
		.blue_n          (hdmi_blue_n),                    //             .blue_n
		.x               (hdmi_x),                         //             .x
		.y               (hdmi_y),                         //             .y
		.horz            (hdmi_horz),                      //             .horz
		.vert            (hdmi_vert),                      //             .vert
		.s_read          (slave_read),                     // avalon_slave.read
		.s_write         (slave_write),                    //             .write
		.s_address       (slave_address),                  //             .address
		.s_writedata     (slave_writedata),                //             .writedata
		.s_burstcount    (slave_burstcount),               //             .burstcount
		.s_byteenable    (slave_byteenable),               //             .byteenable
		.s_waitrequest   (slave_waitrequest),              //             .waitrequest
		.s_readdatavalid (slave_readdatavalid),            //             .readdatavalid
		.s_readdata      (slave_readdata),                 //             .readdata
		.clk_x10         (altpll_0_c0_clk)                 //      clk_x10.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (altpll_0_c1_clk),                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
