


module top_sdram(input clk);

endmodule
