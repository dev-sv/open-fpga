// soc_design_tb.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module soc_design_tb (
	);

	wire         soc_design_inst_clk_bfm_clk_clk;                                        // soc_design_inst_clk_bfm:clk -> [mm_interconnect_0:soc_design_inst_clk_bfm_clk_clk, rst_controller:clk, soc_design_inst:clk_clk, soc_design_inst_hps_0_f2h_axi_slave_bfm:ACLK]
	wire         soc_design_inst_hps_0_f2h_axi_slave_bfm_reset_sink_bfm_clk_bfm_clk_clk; // soc_design_inst_hps_0_f2h_axi_slave_bfm_reset_sink_bfm_clk_bfm:clk -> soc_design_inst_hps_0_f2h_axi_slave_bfm_reset_sink_bfm:clk
	wire         soc_design_inst_hps_io_hps_io_gpio_inst_gpio53;                         // [] -> [soc_design_inst:hps_io_hps_io_gpio_inst_GPIO53, soc_design_inst_hps_io_bfm:sig_hps_io_gpio_inst_GPIO53]
	wire   [0:0] soc_design_inst_memory_bfm_conduit_oct_rzqin;                           // soc_design_inst_memory_bfm:sig_oct_rzqin -> soc_design_inst:memory_oct_rzqin
	wire         soc_design_inst_memory_mem_cas_n;                                       // soc_design_inst:memory_mem_cas_n -> soc_design_inst_memory_bfm:sig_mem_cas_n
	wire         soc_design_inst_memory_mem_reset_n;                                     // soc_design_inst:memory_mem_reset_n -> soc_design_inst_memory_bfm:sig_mem_reset_n
	wire   [2:0] soc_design_inst_memory_mem_ba;                                          // soc_design_inst:memory_mem_ba -> soc_design_inst_memory_bfm:sig_mem_ba
	wire         soc_design_inst_memory_mem_we_n;                                        // soc_design_inst:memory_mem_we_n -> soc_design_inst_memory_bfm:sig_mem_we_n
	wire         soc_design_inst_memory_mem_ck;                                          // soc_design_inst:memory_mem_ck -> soc_design_inst_memory_bfm:sig_mem_ck
	wire   [3:0] soc_design_inst_memory_mem_dm;                                          // soc_design_inst:memory_mem_dm -> soc_design_inst_memory_bfm:sig_mem_dm
	wire   [3:0] soc_design_inst_memory_mem_dqs;                                         // [] -> [soc_design_inst:memory_mem_dqs, soc_design_inst_memory_bfm:sig_mem_dqs]
	wire  [31:0] soc_design_inst_memory_mem_dq;                                          // [] -> [soc_design_inst:memory_mem_dq, soc_design_inst_memory_bfm:sig_mem_dq]
	wire         soc_design_inst_memory_mem_cs_n;                                        // soc_design_inst:memory_mem_cs_n -> soc_design_inst_memory_bfm:sig_mem_cs_n
	wire  [14:0] soc_design_inst_memory_mem_a;                                           // soc_design_inst:memory_mem_a -> soc_design_inst_memory_bfm:sig_mem_a
	wire   [3:0] soc_design_inst_memory_mem_dqs_n;                                       // [] -> [soc_design_inst:memory_mem_dqs_n, soc_design_inst_memory_bfm:sig_mem_dqs_n]
	wire         soc_design_inst_memory_mem_odt;                                         // soc_design_inst:memory_mem_odt -> soc_design_inst_memory_bfm:sig_mem_odt
	wire         soc_design_inst_memory_mem_ras_n;                                       // soc_design_inst:memory_mem_ras_n -> soc_design_inst_memory_bfm:sig_mem_ras_n
	wire         soc_design_inst_memory_mem_ck_n;                                        // soc_design_inst:memory_mem_ck_n -> soc_design_inst_memory_bfm:sig_mem_ck_n
	wire         soc_design_inst_memory_mem_cke;                                         // soc_design_inst:memory_mem_cke -> soc_design_inst_memory_bfm:sig_mem_cke
	wire   [1:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awburst;      // soc_design_inst_hps_0_f2h_axi_slave_bfm:AWBURST -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awburst
	wire   [7:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awuser;       // soc_design_inst_hps_0_f2h_axi_slave_bfm:AWUSER -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awuser
	wire   [3:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arlen;        // soc_design_inst_hps_0_f2h_axi_slave_bfm:ARLEN -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arlen
	wire         soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wready;       // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wready -> soc_design_inst_hps_0_f2h_axi_slave_bfm:WREADY
	wire   [3:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wstrb;        // soc_design_inst_hps_0_f2h_axi_slave_bfm:WSTRB -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wstrb
	wire   [7:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rid;          // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rid -> soc_design_inst_hps_0_f2h_axi_slave_bfm:RID
	wire         soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rready;       // soc_design_inst_hps_0_f2h_axi_slave_bfm:RREADY -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rready
	wire   [3:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awlen;        // soc_design_inst_hps_0_f2h_axi_slave_bfm:AWLEN -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awlen
	wire   [7:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wid;          // soc_design_inst_hps_0_f2h_axi_slave_bfm:WID -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wid
	wire   [3:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arcache;      // soc_design_inst_hps_0_f2h_axi_slave_bfm:ARCACHE -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arcache
	wire         soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wvalid;       // soc_design_inst_hps_0_f2h_axi_slave_bfm:WVALID -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wvalid
	wire  [31:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_araddr;       // soc_design_inst_hps_0_f2h_axi_slave_bfm:ARADDR -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_araddr
	wire   [2:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arprot;       // soc_design_inst_hps_0_f2h_axi_slave_bfm:ARPROT -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arprot
	wire   [2:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awprot;       // soc_design_inst_hps_0_f2h_axi_slave_bfm:AWPROT -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awprot
	wire         soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arvalid;      // soc_design_inst_hps_0_f2h_axi_slave_bfm:ARVALID -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arvalid
	wire  [31:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wdata;        // soc_design_inst_hps_0_f2h_axi_slave_bfm:WDATA -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wdata
	wire   [3:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awcache;      // soc_design_inst_hps_0_f2h_axi_slave_bfm:AWCACHE -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awcache
	wire   [7:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arid;         // soc_design_inst_hps_0_f2h_axi_slave_bfm:ARID -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arid
	wire   [1:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arlock;       // soc_design_inst_hps_0_f2h_axi_slave_bfm:ARLOCK -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arlock
	wire   [1:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awlock;       // soc_design_inst_hps_0_f2h_axi_slave_bfm:AWLOCK -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awlock
	wire  [31:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awaddr;       // soc_design_inst_hps_0_f2h_axi_slave_bfm:AWADDR -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awaddr
	wire         soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arready;      // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arready -> soc_design_inst_hps_0_f2h_axi_slave_bfm:ARREADY
	wire   [1:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_bresp;        // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_bresp -> soc_design_inst_hps_0_f2h_axi_slave_bfm:BRESP
	wire  [31:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rdata;        // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rdata -> soc_design_inst_hps_0_f2h_axi_slave_bfm:RDATA
	wire         soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awready;      // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awready -> soc_design_inst_hps_0_f2h_axi_slave_bfm:AWREADY
	wire   [1:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arburst;      // soc_design_inst_hps_0_f2h_axi_slave_bfm:ARBURST -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arburst
	wire   [2:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arsize;       // soc_design_inst_hps_0_f2h_axi_slave_bfm:ARSIZE -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arsize
	wire         soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rlast;        // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rlast -> soc_design_inst_hps_0_f2h_axi_slave_bfm:RLAST
	wire         soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_bready;       // soc_design_inst_hps_0_f2h_axi_slave_bfm:BREADY -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_bready
	wire         soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wlast;        // soc_design_inst_hps_0_f2h_axi_slave_bfm:WLAST -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wlast
	wire   [1:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rresp;        // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rresp -> soc_design_inst_hps_0_f2h_axi_slave_bfm:RRESP
	wire   [7:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awid;         // soc_design_inst_hps_0_f2h_axi_slave_bfm:AWID -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awid
	wire   [7:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_bid;          // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_bid -> soc_design_inst_hps_0_f2h_axi_slave_bfm:BID
	wire         soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_bvalid;       // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_bvalid -> soc_design_inst_hps_0_f2h_axi_slave_bfm:BVALID
	wire         soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awvalid;      // soc_design_inst_hps_0_f2h_axi_slave_bfm:AWVALID -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awvalid
	wire   [2:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awsize;       // soc_design_inst_hps_0_f2h_axi_slave_bfm:AWSIZE -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awsize
	wire   [7:0] soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_aruser;       // soc_design_inst_hps_0_f2h_axi_slave_bfm:ARUSER -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_aruser
	wire         soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rvalid;       // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rvalid -> soc_design_inst_hps_0_f2h_axi_slave_bfm:RVALID
	wire   [1:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awburst;          // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_awburst -> soc_design_inst:hps_0_f2h_axi_slave_awburst
	wire   [4:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awuser;           // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_awuser -> soc_design_inst:hps_0_f2h_axi_slave_awuser
	wire   [3:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arlen;            // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_arlen -> soc_design_inst:hps_0_f2h_axi_slave_arlen
	wire   [3:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_wstrb;            // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_wstrb -> soc_design_inst:hps_0_f2h_axi_slave_wstrb
	wire         mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_wready;           // soc_design_inst:hps_0_f2h_axi_slave_wready -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_wready
	wire   [7:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_rid;              // soc_design_inst:hps_0_f2h_axi_slave_rid -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_rid
	wire         mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_rready;           // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_rready -> soc_design_inst:hps_0_f2h_axi_slave_rready
	wire   [3:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awlen;            // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_awlen -> soc_design_inst:hps_0_f2h_axi_slave_awlen
	wire   [7:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_wid;              // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_wid -> soc_design_inst:hps_0_f2h_axi_slave_wid
	wire   [3:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arcache;          // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_arcache -> soc_design_inst:hps_0_f2h_axi_slave_arcache
	wire         mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_wvalid;           // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_wvalid -> soc_design_inst:hps_0_f2h_axi_slave_wvalid
	wire  [31:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_araddr;           // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_araddr -> soc_design_inst:hps_0_f2h_axi_slave_araddr
	wire   [2:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arprot;           // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_arprot -> soc_design_inst:hps_0_f2h_axi_slave_arprot
	wire   [2:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awprot;           // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_awprot -> soc_design_inst:hps_0_f2h_axi_slave_awprot
	wire  [31:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_wdata;            // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_wdata -> soc_design_inst:hps_0_f2h_axi_slave_wdata
	wire         mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arvalid;          // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_arvalid -> soc_design_inst:hps_0_f2h_axi_slave_arvalid
	wire   [3:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awcache;          // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_awcache -> soc_design_inst:hps_0_f2h_axi_slave_awcache
	wire   [7:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arid;             // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_arid -> soc_design_inst:hps_0_f2h_axi_slave_arid
	wire   [1:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arlock;           // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_arlock -> soc_design_inst:hps_0_f2h_axi_slave_arlock
	wire   [1:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awlock;           // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_awlock -> soc_design_inst:hps_0_f2h_axi_slave_awlock
	wire  [31:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awaddr;           // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_awaddr -> soc_design_inst:hps_0_f2h_axi_slave_awaddr
	wire   [1:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_bresp;            // soc_design_inst:hps_0_f2h_axi_slave_bresp -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bresp
	wire         mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arready;          // soc_design_inst:hps_0_f2h_axi_slave_arready -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_arready
	wire  [31:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_rdata;            // soc_design_inst:hps_0_f2h_axi_slave_rdata -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_rdata
	wire         mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awready;          // soc_design_inst:hps_0_f2h_axi_slave_awready -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_awready
	wire   [1:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arburst;          // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_arburst -> soc_design_inst:hps_0_f2h_axi_slave_arburst
	wire   [2:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arsize;           // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_arsize -> soc_design_inst:hps_0_f2h_axi_slave_arsize
	wire         mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_bready;           // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bready -> soc_design_inst:hps_0_f2h_axi_slave_bready
	wire         mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_rlast;            // soc_design_inst:hps_0_f2h_axi_slave_rlast -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_rlast
	wire         mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_wlast;            // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_wlast -> soc_design_inst:hps_0_f2h_axi_slave_wlast
	wire   [1:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_rresp;            // soc_design_inst:hps_0_f2h_axi_slave_rresp -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_rresp
	wire   [7:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awid;             // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_awid -> soc_design_inst:hps_0_f2h_axi_slave_awid
	wire   [7:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_bid;              // soc_design_inst:hps_0_f2h_axi_slave_bid -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bid
	wire         mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_bvalid;           // soc_design_inst:hps_0_f2h_axi_slave_bvalid -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bvalid
	wire   [2:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awsize;           // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_awsize -> soc_design_inst:hps_0_f2h_axi_slave_awsize
	wire         mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awvalid;          // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_awvalid -> soc_design_inst:hps_0_f2h_axi_slave_awvalid
	wire   [4:0] mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_aruser;           // mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_aruser -> soc_design_inst:hps_0_f2h_axi_slave_aruser
	wire         mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_rvalid;           // soc_design_inst:hps_0_f2h_axi_slave_rvalid -> mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_rvalid
	wire         rst_controller_reset_out_reset;                                         // rst_controller:reset_out -> [mm_interconnect_0:soc_design_inst_hps_0_f2h_axi_slave_bfm_reset_sink_reset_bridge_in_reset_reset, soc_design_inst_hps_0_f2h_axi_slave_bfm:ARESETn]
	wire         soc_design_inst_hps_0_f2h_axi_slave_bfm_reset_sink_bfm_reset_reset;     // soc_design_inst_hps_0_f2h_axi_slave_bfm_reset_sink_bfm:reset -> rst_controller:reset_in0

	soc_design soc_design_inst (
		.clk_clk                        (soc_design_inst_clk_bfm_clk_clk),                               //                 clk.clk
		.hps_0_f2h_axi_slave_awid       (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awid),    // hps_0_f2h_axi_slave.awid
		.hps_0_f2h_axi_slave_awaddr     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awaddr),  //                    .awaddr
		.hps_0_f2h_axi_slave_awlen      (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awlen),   //                    .awlen
		.hps_0_f2h_axi_slave_awsize     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awsize),  //                    .awsize
		.hps_0_f2h_axi_slave_awburst    (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awburst), //                    .awburst
		.hps_0_f2h_axi_slave_awlock     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awlock),  //                    .awlock
		.hps_0_f2h_axi_slave_awcache    (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awcache), //                    .awcache
		.hps_0_f2h_axi_slave_awprot     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awprot),  //                    .awprot
		.hps_0_f2h_axi_slave_awvalid    (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awvalid), //                    .awvalid
		.hps_0_f2h_axi_slave_awready    (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awready), //                    .awready
		.hps_0_f2h_axi_slave_awuser     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awuser),  //                    .awuser
		.hps_0_f2h_axi_slave_wid        (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_wid),     //                    .wid
		.hps_0_f2h_axi_slave_wdata      (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_wdata),   //                    .wdata
		.hps_0_f2h_axi_slave_wstrb      (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_wstrb),   //                    .wstrb
		.hps_0_f2h_axi_slave_wlast      (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_wlast),   //                    .wlast
		.hps_0_f2h_axi_slave_wvalid     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_wvalid),  //                    .wvalid
		.hps_0_f2h_axi_slave_wready     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_wready),  //                    .wready
		.hps_0_f2h_axi_slave_bid        (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_bid),     //                    .bid
		.hps_0_f2h_axi_slave_bresp      (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_bresp),   //                    .bresp
		.hps_0_f2h_axi_slave_bvalid     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_bvalid),  //                    .bvalid
		.hps_0_f2h_axi_slave_bready     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_bready),  //                    .bready
		.hps_0_f2h_axi_slave_arid       (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arid),    //                    .arid
		.hps_0_f2h_axi_slave_araddr     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_araddr),  //                    .araddr
		.hps_0_f2h_axi_slave_arlen      (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arlen),   //                    .arlen
		.hps_0_f2h_axi_slave_arsize     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arsize),  //                    .arsize
		.hps_0_f2h_axi_slave_arburst    (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arburst), //                    .arburst
		.hps_0_f2h_axi_slave_arlock     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arlock),  //                    .arlock
		.hps_0_f2h_axi_slave_arcache    (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arcache), //                    .arcache
		.hps_0_f2h_axi_slave_arprot     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arprot),  //                    .arprot
		.hps_0_f2h_axi_slave_arvalid    (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arvalid), //                    .arvalid
		.hps_0_f2h_axi_slave_arready    (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arready), //                    .arready
		.hps_0_f2h_axi_slave_aruser     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_aruser),  //                    .aruser
		.hps_0_f2h_axi_slave_rid        (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_rid),     //                    .rid
		.hps_0_f2h_axi_slave_rdata      (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_rdata),   //                    .rdata
		.hps_0_f2h_axi_slave_rresp      (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_rresp),   //                    .rresp
		.hps_0_f2h_axi_slave_rlast      (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_rlast),   //                    .rlast
		.hps_0_f2h_axi_slave_rvalid     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_rvalid),  //                    .rvalid
		.hps_0_f2h_axi_slave_rready     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_rready),  //                    .rready
		.hps_io_hps_io_gpio_inst_GPIO53 (soc_design_inst_hps_io_hps_io_gpio_inst_gpio53),                //              hps_io.hps_io_gpio_inst_GPIO53
		.memory_mem_a                   (soc_design_inst_memory_mem_a),                                  //              memory.mem_a
		.memory_mem_ba                  (soc_design_inst_memory_mem_ba),                                 //                    .mem_ba
		.memory_mem_ck                  (soc_design_inst_memory_mem_ck),                                 //                    .mem_ck
		.memory_mem_ck_n                (soc_design_inst_memory_mem_ck_n),                               //                    .mem_ck_n
		.memory_mem_cke                 (soc_design_inst_memory_mem_cke),                                //                    .mem_cke
		.memory_mem_cs_n                (soc_design_inst_memory_mem_cs_n),                               //                    .mem_cs_n
		.memory_mem_ras_n               (soc_design_inst_memory_mem_ras_n),                              //                    .mem_ras_n
		.memory_mem_cas_n               (soc_design_inst_memory_mem_cas_n),                              //                    .mem_cas_n
		.memory_mem_we_n                (soc_design_inst_memory_mem_we_n),                               //                    .mem_we_n
		.memory_mem_reset_n             (soc_design_inst_memory_mem_reset_n),                            //                    .mem_reset_n
		.memory_mem_dq                  (soc_design_inst_memory_mem_dq),                                 //                    .mem_dq
		.memory_mem_dqs                 (soc_design_inst_memory_mem_dqs),                                //                    .mem_dqs
		.memory_mem_dqs_n               (soc_design_inst_memory_mem_dqs_n),                              //                    .mem_dqs_n
		.memory_mem_odt                 (soc_design_inst_memory_mem_odt),                                //                    .mem_odt
		.memory_mem_dm                  (soc_design_inst_memory_mem_dm),                                 //                    .mem_dm
		.memory_oct_rzqin               (soc_design_inst_memory_bfm_conduit_oct_rzqin)                   //                    .oct_rzqin
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) soc_design_inst_clk_bfm (
		.clk (soc_design_inst_clk_bfm_clk_clk)  // clk.clk
	);

	mgc_axi_master #(
		.AXI_ADDRESS_WIDTH           (32),
		.AXI_RDATA_WIDTH             (32),
		.AXI_WDATA_WIDTH             (32),
		.AXI_ID_WIDTH                (8),
		.index                       (0),
		.READ_ISSUING_CAPABILITY     (16),
		.WRITE_ISSUING_CAPABILITY    (16),
		.COMBINED_ISSUING_CAPABILITY (16)
	) soc_design_inst_hps_0_f2h_axi_slave_bfm (
		.AWVALID (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awvalid), // altera_axi_master.awvalid
		.AWLEN   (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awlen),   //                  .awlen
		.AWSIZE  (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awsize),  //                  .awsize
		.AWBURST (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awburst), //                  .awburst
		.AWLOCK  (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awlock),  //                  .awlock
		.AWCACHE (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awcache), //                  .awcache
		.AWPROT  (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awprot),  //                  .awprot
		.AWREADY (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awready), //                  .awready
		.AWUSER  (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awuser),  //                  .awuser
		.ARVALID (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arvalid), //                  .arvalid
		.ARLEN   (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arlen),   //                  .arlen
		.ARSIZE  (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arsize),  //                  .arsize
		.ARBURST (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arburst), //                  .arburst
		.ARLOCK  (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arlock),  //                  .arlock
		.ARCACHE (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arcache), //                  .arcache
		.ARPROT  (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arprot),  //                  .arprot
		.ARREADY (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arready), //                  .arready
		.ARUSER  (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_aruser),  //                  .aruser
		.RVALID  (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rvalid),  //                  .rvalid
		.RLAST   (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rlast),   //                  .rlast
		.RRESP   (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rresp),   //                  .rresp
		.RREADY  (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rready),  //                  .rready
		.WVALID  (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wvalid),  //                  .wvalid
		.WLAST   (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wlast),   //                  .wlast
		.WREADY  (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wready),  //                  .wready
		.BVALID  (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_bvalid),  //                  .bvalid
		.BRESP   (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_bresp),   //                  .bresp
		.BREADY  (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_bready),  //                  .bready
		.AWADDR  (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awaddr),  //                  .awaddr
		.AWID    (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awid),    //                  .awid
		.ARADDR  (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_araddr),  //                  .araddr
		.ARID    (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arid),    //                  .arid
		.RDATA   (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rdata),   //                  .rdata
		.RID     (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rid),     //                  .rid
		.WDATA   (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wdata),   //                  .wdata
		.WSTRB   (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wstrb),   //                  .wstrb
		.WID     (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wid),     //                  .wid
		.BID     (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_bid),     //                  .bid
		.ACLK    (soc_design_inst_clk_bfm_clk_clk),                                   //        clock_sink.clk
		.ARESETn (~rst_controller_reset_out_reset)                                    //        reset_sink.reset_n
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) soc_design_inst_hps_0_f2h_axi_slave_bfm_reset_sink_bfm (
		.reset (soc_design_inst_hps_0_f2h_axi_slave_bfm_reset_sink_bfm_reset_reset),     // reset.reset_n
		.clk   (soc_design_inst_hps_0_f2h_axi_slave_bfm_reset_sink_bfm_clk_bfm_clk_clk)  //   clk.clk
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) soc_design_inst_hps_0_f2h_axi_slave_bfm_reset_sink_bfm_clk_bfm (
		.clk (soc_design_inst_hps_0_f2h_axi_slave_bfm_reset_sink_bfm_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm soc_design_inst_hps_io_bfm (
		.sig_hps_io_gpio_inst_GPIO53 (soc_design_inst_hps_io_hps_io_gpio_inst_gpio53)  // conduit.hps_io_gpio_inst_GPIO53
	);

	altera_conduit_bfm_0002 soc_design_inst_memory_bfm (
		.sig_mem_a       (soc_design_inst_memory_mem_a),                 // conduit.mem_a
		.sig_mem_ba      (soc_design_inst_memory_mem_ba),                //        .mem_ba
		.sig_mem_cas_n   (soc_design_inst_memory_mem_cas_n),             //        .mem_cas_n
		.sig_mem_ck      (soc_design_inst_memory_mem_ck),                //        .mem_ck
		.sig_mem_ck_n    (soc_design_inst_memory_mem_ck_n),              //        .mem_ck_n
		.sig_mem_cke     (soc_design_inst_memory_mem_cke),               //        .mem_cke
		.sig_mem_cs_n    (soc_design_inst_memory_mem_cs_n),              //        .mem_cs_n
		.sig_mem_dm      (soc_design_inst_memory_mem_dm),                //        .mem_dm
		.sig_mem_dq      (soc_design_inst_memory_mem_dq),                //        .mem_dq
		.sig_mem_dqs     (soc_design_inst_memory_mem_dqs),               //        .mem_dqs
		.sig_mem_dqs_n   (soc_design_inst_memory_mem_dqs_n),             //        .mem_dqs_n
		.sig_mem_odt     (soc_design_inst_memory_mem_odt),               //        .mem_odt
		.sig_mem_ras_n   (soc_design_inst_memory_mem_ras_n),             //        .mem_ras_n
		.sig_mem_reset_n (soc_design_inst_memory_mem_reset_n),           //        .mem_reset_n
		.sig_mem_we_n    (soc_design_inst_memory_mem_we_n),              //        .mem_we_n
		.sig_oct_rzqin   (soc_design_inst_memory_bfm_conduit_oct_rzqin)  //        .oct_rzqin
	);

	altera_mm_interconnect mm_interconnect_0 (
		.soc_design_inst_hps_0_f2h_axi_slave_awid                                       (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awid),        //                                      soc_design_inst_hps_0_f2h_axi_slave.awid
		.soc_design_inst_hps_0_f2h_axi_slave_awaddr                                     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awaddr),      //                                                                         .awaddr
		.soc_design_inst_hps_0_f2h_axi_slave_awlen                                      (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awlen),       //                                                                         .awlen
		.soc_design_inst_hps_0_f2h_axi_slave_awsize                                     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awsize),      //                                                                         .awsize
		.soc_design_inst_hps_0_f2h_axi_slave_awburst                                    (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awburst),     //                                                                         .awburst
		.soc_design_inst_hps_0_f2h_axi_slave_awlock                                     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awlock),      //                                                                         .awlock
		.soc_design_inst_hps_0_f2h_axi_slave_awcache                                    (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awcache),     //                                                                         .awcache
		.soc_design_inst_hps_0_f2h_axi_slave_awprot                                     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awprot),      //                                                                         .awprot
		.soc_design_inst_hps_0_f2h_axi_slave_awuser                                     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awuser),      //                                                                         .awuser
		.soc_design_inst_hps_0_f2h_axi_slave_awvalid                                    (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awvalid),     //                                                                         .awvalid
		.soc_design_inst_hps_0_f2h_axi_slave_awready                                    (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_awready),     //                                                                         .awready
		.soc_design_inst_hps_0_f2h_axi_slave_wid                                        (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_wid),         //                                                                         .wid
		.soc_design_inst_hps_0_f2h_axi_slave_wdata                                      (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_wdata),       //                                                                         .wdata
		.soc_design_inst_hps_0_f2h_axi_slave_wstrb                                      (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_wstrb),       //                                                                         .wstrb
		.soc_design_inst_hps_0_f2h_axi_slave_wlast                                      (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_wlast),       //                                                                         .wlast
		.soc_design_inst_hps_0_f2h_axi_slave_wvalid                                     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_wvalid),      //                                                                         .wvalid
		.soc_design_inst_hps_0_f2h_axi_slave_wready                                     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_wready),      //                                                                         .wready
		.soc_design_inst_hps_0_f2h_axi_slave_bid                                        (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_bid),         //                                                                         .bid
		.soc_design_inst_hps_0_f2h_axi_slave_bresp                                      (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_bresp),       //                                                                         .bresp
		.soc_design_inst_hps_0_f2h_axi_slave_bvalid                                     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_bvalid),      //                                                                         .bvalid
		.soc_design_inst_hps_0_f2h_axi_slave_bready                                     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_bready),      //                                                                         .bready
		.soc_design_inst_hps_0_f2h_axi_slave_arid                                       (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arid),        //                                                                         .arid
		.soc_design_inst_hps_0_f2h_axi_slave_araddr                                     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_araddr),      //                                                                         .araddr
		.soc_design_inst_hps_0_f2h_axi_slave_arlen                                      (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arlen),       //                                                                         .arlen
		.soc_design_inst_hps_0_f2h_axi_slave_arsize                                     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arsize),      //                                                                         .arsize
		.soc_design_inst_hps_0_f2h_axi_slave_arburst                                    (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arburst),     //                                                                         .arburst
		.soc_design_inst_hps_0_f2h_axi_slave_arlock                                     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arlock),      //                                                                         .arlock
		.soc_design_inst_hps_0_f2h_axi_slave_arcache                                    (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arcache),     //                                                                         .arcache
		.soc_design_inst_hps_0_f2h_axi_slave_arprot                                     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arprot),      //                                                                         .arprot
		.soc_design_inst_hps_0_f2h_axi_slave_aruser                                     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_aruser),      //                                                                         .aruser
		.soc_design_inst_hps_0_f2h_axi_slave_arvalid                                    (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arvalid),     //                                                                         .arvalid
		.soc_design_inst_hps_0_f2h_axi_slave_arready                                    (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_arready),     //                                                                         .arready
		.soc_design_inst_hps_0_f2h_axi_slave_rid                                        (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_rid),         //                                                                         .rid
		.soc_design_inst_hps_0_f2h_axi_slave_rdata                                      (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_rdata),       //                                                                         .rdata
		.soc_design_inst_hps_0_f2h_axi_slave_rresp                                      (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_rresp),       //                                                                         .rresp
		.soc_design_inst_hps_0_f2h_axi_slave_rlast                                      (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_rlast),       //                                                                         .rlast
		.soc_design_inst_hps_0_f2h_axi_slave_rvalid                                     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_rvalid),      //                                                                         .rvalid
		.soc_design_inst_hps_0_f2h_axi_slave_rready                                     (mm_interconnect_0_soc_design_inst_hps_0_f2h_axi_slave_rready),      //                                                                         .rready
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awid                 (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awid),    //                soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master.awid
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awaddr               (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awaddr),  //                                                                         .awaddr
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awlen                (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awlen),   //                                                                         .awlen
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awsize               (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awsize),  //                                                                         .awsize
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awburst              (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awburst), //                                                                         .awburst
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awlock               (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awlock),  //                                                                         .awlock
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awcache              (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awcache), //                                                                         .awcache
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awprot               (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awprot),  //                                                                         .awprot
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awuser               (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awuser),  //                                                                         .awuser
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awvalid              (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awvalid), //                                                                         .awvalid
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awready              (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_awready), //                                                                         .awready
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wid                  (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wid),     //                                                                         .wid
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wdata                (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wdata),   //                                                                         .wdata
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wstrb                (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wstrb),   //                                                                         .wstrb
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wlast                (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wlast),   //                                                                         .wlast
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wvalid               (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wvalid),  //                                                                         .wvalid
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wready               (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_wready),  //                                                                         .wready
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_bid                  (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_bid),     //                                                                         .bid
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_bresp                (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_bresp),   //                                                                         .bresp
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_bvalid               (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_bvalid),  //                                                                         .bvalid
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_bready               (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_bready),  //                                                                         .bready
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arid                 (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arid),    //                                                                         .arid
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_araddr               (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_araddr),  //                                                                         .araddr
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arlen                (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arlen),   //                                                                         .arlen
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arsize               (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arsize),  //                                                                         .arsize
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arburst              (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arburst), //                                                                         .arburst
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arlock               (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arlock),  //                                                                         .arlock
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arcache              (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arcache), //                                                                         .arcache
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arprot               (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arprot),  //                                                                         .arprot
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_aruser               (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_aruser),  //                                                                         .aruser
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arvalid              (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arvalid), //                                                                         .arvalid
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arready              (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_arready), //                                                                         .arready
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rid                  (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rid),     //                                                                         .rid
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rdata                (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rdata),   //                                                                         .rdata
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rresp                (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rresp),   //                                                                         .rresp
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rlast                (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rlast),   //                                                                         .rlast
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rvalid               (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rvalid),  //                                                                         .rvalid
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rready               (soc_design_inst_hps_0_f2h_axi_slave_bfm_altera_axi_master_rready),  //                                                                         .rready
		.soc_design_inst_clk_bfm_clk_clk                                                (soc_design_inst_clk_bfm_clk_clk),                                   //                                              soc_design_inst_clk_bfm_clk.clk
		.soc_design_inst_hps_0_f2h_axi_slave_bfm_reset_sink_reset_bridge_in_reset_reset (rst_controller_reset_out_reset)                                     // soc_design_inst_hps_0_f2h_axi_slave_bfm_reset_sink_reset_bridge_in_reset.reset
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~soc_design_inst_hps_0_f2h_axi_slave_bfm_reset_sink_bfm_reset_reset), // reset_in0.reset
		.clk            (soc_design_inst_clk_bfm_clk_clk),                                     //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),                                      // reset_out.reset
		.reset_req      (),                                                                    // (terminated)
		.reset_req_in0  (1'b0),                                                                // (terminated)
		.reset_in1      (1'b0),                                                                // (terminated)
		.reset_req_in1  (1'b0),                                                                // (terminated)
		.reset_in2      (1'b0),                                                                // (terminated)
		.reset_req_in2  (1'b0),                                                                // (terminated)
		.reset_in3      (1'b0),                                                                // (terminated)
		.reset_req_in3  (1'b0),                                                                // (terminated)
		.reset_in4      (1'b0),                                                                // (terminated)
		.reset_req_in4  (1'b0),                                                                // (terminated)
		.reset_in5      (1'b0),                                                                // (terminated)
		.reset_req_in5  (1'b0),                                                                // (terminated)
		.reset_in6      (1'b0),                                                                // (terminated)
		.reset_req_in6  (1'b0),                                                                // (terminated)
		.reset_in7      (1'b0),                                                                // (terminated)
		.reset_req_in7  (1'b0),                                                                // (terminated)
		.reset_in8      (1'b0),                                                                // (terminated)
		.reset_req_in8  (1'b0),                                                                // (terminated)
		.reset_in9      (1'b0),                                                                // (terminated)
		.reset_req_in9  (1'b0),                                                                // (terminated)
		.reset_in10     (1'b0),                                                                // (terminated)
		.reset_req_in10 (1'b0),                                                                // (terminated)
		.reset_in11     (1'b0),                                                                // (terminated)
		.reset_req_in11 (1'b0),                                                                // (terminated)
		.reset_in12     (1'b0),                                                                // (terminated)
		.reset_req_in12 (1'b0),                                                                // (terminated)
		.reset_in13     (1'b0),                                                                // (terminated)
		.reset_req_in13 (1'b0),                                                                // (terminated)
		.reset_in14     (1'b0),                                                                // (terminated)
		.reset_req_in14 (1'b0),                                                                // (terminated)
		.reset_in15     (1'b0),                                                                // (terminated)
		.reset_req_in15 (1'b0)                                                                 // (terminated)
	);

endmodule
