// soc_design.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module soc_design (
		input  wire        clk_clk,            //    clk.clk
		output wire [12:0] memory_mem_a,       // memory.mem_a
		output wire [2:0]  memory_mem_ba,      //       .mem_ba
		output wire        memory_mem_ck,      //       .mem_ck
		output wire        memory_mem_ck_n,    //       .mem_ck_n
		output wire        memory_mem_cke,     //       .mem_cke
		output wire        memory_mem_cs_n,    //       .mem_cs_n
		output wire        memory_mem_ras_n,   //       .mem_ras_n
		output wire        memory_mem_cas_n,   //       .mem_cas_n
		output wire        memory_mem_we_n,    //       .mem_we_n
		output wire        memory_mem_reset_n, //       .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,      //       .mem_dq
		inout  wire        memory_mem_dqs,     //       .mem_dqs
		inout  wire        memory_mem_dqs_n,   //       .mem_dqs_n
		output wire        memory_mem_odt,     //       .mem_odt
		output wire        memory_mem_dm,      //       .mem_dm
		input  wire        memory_oct_rzqin,   //       .oct_rzqin
		input  wire        reset_reset_n       //  reset.reset_n
	);

	soc_design_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (0)
	) hps_0 (
		.mem_a                    (memory_mem_a),       //           memory.mem_a
		.mem_ba                   (memory_mem_ba),      //                 .mem_ba
		.mem_ck                   (memory_mem_ck),      //                 .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),    //                 .mem_ck_n
		.mem_cke                  (memory_mem_cke),     //                 .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),    //                 .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),   //                 .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),   //                 .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),    //                 .mem_we_n
		.mem_reset_n              (memory_mem_reset_n), //                 .mem_reset_n
		.mem_dq                   (memory_mem_dq),      //                 .mem_dq
		.mem_dqs                  (memory_mem_dqs),     //                 .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),   //                 .mem_dqs_n
		.mem_odt                  (memory_mem_odt),     //                 .mem_odt
		.mem_dm                   (memory_mem_dm),      //                 .mem_dm
		.oct_rzqin                (memory_oct_rzqin),   //                 .oct_rzqin
		.h2f_rst_n                (),                   //        h2f_reset.reset_n
		.f2h_sdram0_clk           (clk_clk),            // f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS       (),                   //  f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT    (),                   //                 .burstcount
		.f2h_sdram0_WAITREQUEST   (),                   //                 .waitrequest
		.f2h_sdram0_READDATA      (),                   //                 .readdata
		.f2h_sdram0_READDATAVALID (),                   //                 .readdatavalid
		.f2h_sdram0_READ          ()                    //                 .read
	);

endmodule
