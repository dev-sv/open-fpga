


module button(input bit clk);





endmodule: button