// avl_if.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module avl_if (
		input  wire        aclk_aclk,         //  aclk.aclk
		output wire        adc_waitrequest,   //   adc.waitrequest
		output wire [15:0] adc_readdata,      //      .readdata
		output wire        adc_readdatavalid, //      .readdatavalid
		input  wire [0:0]  adc_burstcount,    //      .burstcount
		input  wire [15:0] adc_writedata,     //      .writedata
		input  wire [9:0]  adc_address,       //      .address
		input  wire        adc_write,         //      .write
		input  wire        adc_read,          //      .read
		input  wire [1:0]  adc_byteenable,    //      .byteenable
		input  wire        adc_debugaccess,   //      .debugaccess
		input  wire        clk_clk,           //   clk.clk
		input  wire        reset_reset_n      // reset.reset_n
	);

	wire         mm_bridge_0_m0_waitrequest;                                 // mm_interconnect_0:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	wire  [15:0] mm_bridge_0_m0_readdata;                                    // mm_interconnect_0:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	wire         mm_bridge_0_m0_debugaccess;                                 // mm_bridge_0:m0_debugaccess -> mm_interconnect_0:mm_bridge_0_m0_debugaccess
	wire   [9:0] mm_bridge_0_m0_address;                                     // mm_bridge_0:m0_address -> mm_interconnect_0:mm_bridge_0_m0_address
	wire         mm_bridge_0_m0_read;                                        // mm_bridge_0:m0_read -> mm_interconnect_0:mm_bridge_0_m0_read
	wire   [1:0] mm_bridge_0_m0_byteenable;                                  // mm_bridge_0:m0_byteenable -> mm_interconnect_0:mm_bridge_0_m0_byteenable
	wire         mm_bridge_0_m0_readdatavalid;                               // mm_interconnect_0:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	wire  [15:0] mm_bridge_0_m0_writedata;                                   // mm_bridge_0:m0_writedata -> mm_interconnect_0:mm_bridge_0_m0_writedata
	wire         mm_bridge_0_m0_write;                                       // mm_bridge_0:m0_write -> mm_interconnect_0:mm_bridge_0_m0_write
	wire   [0:0] mm_bridge_0_m0_burstcount;                                  // mm_bridge_0:m0_burstcount -> mm_interconnect_0:mm_bridge_0_m0_burstcount
	wire  [15:0] mm_interconnect_0_adc_max10_0_avalon_slave_0_readdata;      // adc_max10_0:readdata -> mm_interconnect_0:adc_max10_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_adc_max10_0_avalon_slave_0_waitrequest;   // adc_max10_0:waitrequest -> mm_interconnect_0:adc_max10_0_avalon_slave_0_waitrequest
	wire   [9:0] mm_interconnect_0_adc_max10_0_avalon_slave_0_address;       // mm_interconnect_0:adc_max10_0_avalon_slave_0_address -> adc_max10_0:address
	wire         mm_interconnect_0_adc_max10_0_avalon_slave_0_read;          // mm_interconnect_0:adc_max10_0_avalon_slave_0_read -> adc_max10_0:read
	wire         mm_interconnect_0_adc_max10_0_avalon_slave_0_readdatavalid; // adc_max10_0:readdatavalid -> mm_interconnect_0:adc_max10_0_avalon_slave_0_readdatavalid
	wire         mm_interconnect_0_adc_max10_0_avalon_slave_0_write;         // mm_interconnect_0:adc_max10_0_avalon_slave_0_write -> adc_max10_0:write
	wire  [15:0] mm_interconnect_0_adc_max10_0_avalon_slave_0_writedata;     // mm_interconnect_0:adc_max10_0_avalon_slave_0_writedata -> adc_max10_0:writedata
	wire   [0:0] mm_interconnect_0_adc_max10_0_avalon_slave_0_burstcount;    // mm_interconnect_0:adc_max10_0_avalon_slave_0_burstcount -> adc_max10_0:burstcount
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [adc_max10_0:reset, mm_bridge_0:reset, mm_interconnect_0:mm_bridge_0_reset_reset_bridge_in_reset_reset]

	adc adc_max10_0 (
		.clk           (clk_clk),                                                    //          clock.clk
		.reset         (rst_controller_reset_out_reset),                             //          reset.reset
		.write         (mm_interconnect_0_adc_max10_0_avalon_slave_0_write),         // avalon_slave_0.write
		.read          (mm_interconnect_0_adc_max10_0_avalon_slave_0_read),          //               .read
		.address       (mm_interconnect_0_adc_max10_0_avalon_slave_0_address),       //               .address
		.writedata     (mm_interconnect_0_adc_max10_0_avalon_slave_0_writedata),     //               .writedata
		.readdata      (mm_interconnect_0_adc_max10_0_avalon_slave_0_readdata),      //               .readdata
		.readdatavalid (mm_interconnect_0_adc_max10_0_avalon_slave_0_readdatavalid), //               .readdatavalid
		.burstcount    (mm_interconnect_0_adc_max10_0_avalon_slave_0_burstcount),    //               .burstcount
		.waitrequest   (mm_interconnect_0_adc_max10_0_avalon_slave_0_waitrequest),   //               .waitrequest
		.aclk          (aclk_aclk)                                                   //           aclk.aclk
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (16),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (10),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_0 (
		.clk              (clk_clk),                        //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (adc_waitrequest),                //    s0.waitrequest
		.s0_readdata      (adc_readdata),                   //      .readdata
		.s0_readdatavalid (adc_readdatavalid),              //      .readdatavalid
		.s0_burstcount    (adc_burstcount),                 //      .burstcount
		.s0_writedata     (adc_writedata),                  //      .writedata
		.s0_address       (adc_address),                    //      .address
		.s0_write         (adc_write),                      //      .write
		.s0_read          (adc_read),                       //      .read
		.s0_byteenable    (adc_byteenable),                 //      .byteenable
		.s0_debugaccess   (adc_debugaccess),                //      .debugaccess
		.m0_waitrequest   (mm_bridge_0_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_0_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_0_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_0_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_0_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_0_m0_address),         //      .address
		.m0_write         (mm_bridge_0_m0_write),           //      .write
		.m0_read          (mm_bridge_0_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_0_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_0_m0_debugaccess),     //      .debugaccess
		.s0_response      (),                               // (terminated)
		.m0_response      (2'b00)                           // (terminated)
	);

	avl_if_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                 (clk_clk),                                                    //                               clk_0_clk.clk
		.mm_bridge_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                             // mm_bridge_0_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_m0_address                        (mm_bridge_0_m0_address),                                     //                          mm_bridge_0_m0.address
		.mm_bridge_0_m0_waitrequest                    (mm_bridge_0_m0_waitrequest),                                 //                                        .waitrequest
		.mm_bridge_0_m0_burstcount                     (mm_bridge_0_m0_burstcount),                                  //                                        .burstcount
		.mm_bridge_0_m0_byteenable                     (mm_bridge_0_m0_byteenable),                                  //                                        .byteenable
		.mm_bridge_0_m0_read                           (mm_bridge_0_m0_read),                                        //                                        .read
		.mm_bridge_0_m0_readdata                       (mm_bridge_0_m0_readdata),                                    //                                        .readdata
		.mm_bridge_0_m0_readdatavalid                  (mm_bridge_0_m0_readdatavalid),                               //                                        .readdatavalid
		.mm_bridge_0_m0_write                          (mm_bridge_0_m0_write),                                       //                                        .write
		.mm_bridge_0_m0_writedata                      (mm_bridge_0_m0_writedata),                                   //                                        .writedata
		.mm_bridge_0_m0_debugaccess                    (mm_bridge_0_m0_debugaccess),                                 //                                        .debugaccess
		.adc_max10_0_avalon_slave_0_address            (mm_interconnect_0_adc_max10_0_avalon_slave_0_address),       //              adc_max10_0_avalon_slave_0.address
		.adc_max10_0_avalon_slave_0_write              (mm_interconnect_0_adc_max10_0_avalon_slave_0_write),         //                                        .write
		.adc_max10_0_avalon_slave_0_read               (mm_interconnect_0_adc_max10_0_avalon_slave_0_read),          //                                        .read
		.adc_max10_0_avalon_slave_0_readdata           (mm_interconnect_0_adc_max10_0_avalon_slave_0_readdata),      //                                        .readdata
		.adc_max10_0_avalon_slave_0_writedata          (mm_interconnect_0_adc_max10_0_avalon_slave_0_writedata),     //                                        .writedata
		.adc_max10_0_avalon_slave_0_burstcount         (mm_interconnect_0_adc_max10_0_avalon_slave_0_burstcount),    //                                        .burstcount
		.adc_max10_0_avalon_slave_0_readdatavalid      (mm_interconnect_0_adc_max10_0_avalon_slave_0_readdatavalid), //                                        .readdatavalid
		.adc_max10_0_avalon_slave_0_waitrequest        (mm_interconnect_0_adc_max10_0_avalon_slave_0_waitrequest)    //                                        .waitrequest
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
