
module adc_qsys (
	aclk_clk,
	clk_clk,
	reset_reset_n);	

	input		aclk_clk;
	input		clk_clk;
	input		reset_reset_n;
endmodule
