


module tb_top(input clk);


endmodule
