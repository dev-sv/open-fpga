


module adc_ip(input clk);

endmodule
