// hdmi_qsys.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module hdmi_qsys (
		input  wire        clk_clk,        //     clk.clk
		input  wire        clk_x10_clk,    // clk_x10.clk
		output wire        hdmi_clk_mm,    //    hdmi.clk_mm
		output wire        hdmi_clk_pix_p, //        .clk_pix_p
		output wire        hdmi_clk_pix_n, //        .clk_pix_n
		output wire        hdmi_red_p,     //        .red_p
		output wire        hdmi_red_n,     //        .red_n
		output wire        hdmi_green_p,   //        .green_p
		output wire        hdmi_green_n,   //        .green_n
		output wire        hdmi_blue_p,    //        .blue_p
		output wire        hdmi_blue_n,    //        .blue_n
		output wire [10:0] hdmi_x,         //        .x
		output wire [10:0] hdmi_y,         //        .y
		output wire [10:0] hdmi_horz,      //        .horz
		output wire [10:0] hdmi_vert,      //        .vert
		input  wire        reset_reset_n   //   reset.reset_n
	);

	wire  [31:0] master_bfm_m0_readdata;                               // mm_interconnect_0:master_bfm_m0_readdata -> master_bfm:avm_readdata
	wire         master_bfm_m0_waitrequest;                            // mm_interconnect_0:master_bfm_m0_waitrequest -> master_bfm:avm_waitrequest
	wire  [31:0] master_bfm_m0_address;                                // master_bfm:avm_address -> mm_interconnect_0:master_bfm_m0_address
	wire         master_bfm_m0_read;                                   // master_bfm:avm_read -> mm_interconnect_0:master_bfm_m0_read
	wire   [3:0] master_bfm_m0_byteenable;                             // master_bfm:avm_byteenable -> mm_interconnect_0:master_bfm_m0_byteenable
	wire         master_bfm_m0_readdatavalid;                          // mm_interconnect_0:master_bfm_m0_readdatavalid -> master_bfm:avm_readdatavalid
	wire  [31:0] master_bfm_m0_writedata;                              // master_bfm:avm_writedata -> mm_interconnect_0:master_bfm_m0_writedata
	wire         master_bfm_m0_write;                                  // master_bfm:avm_write -> mm_interconnect_0:master_bfm_m0_write
	wire   [0:0] master_bfm_m0_burstcount;                             // master_bfm:avm_burstcount -> mm_interconnect_0:master_bfm_m0_burstcount
	wire  [31:0] mm_interconnect_0_hdmi_mm_avalon_slave_readdata;      // hdmi_mm:s_readdata -> mm_interconnect_0:hdmi_mm_avalon_slave_readdata
	wire         mm_interconnect_0_hdmi_mm_avalon_slave_waitrequest;   // hdmi_mm:s_waitrequest -> mm_interconnect_0:hdmi_mm_avalon_slave_waitrequest
	wire   [9:0] mm_interconnect_0_hdmi_mm_avalon_slave_address;       // mm_interconnect_0:hdmi_mm_avalon_slave_address -> hdmi_mm:s_address
	wire         mm_interconnect_0_hdmi_mm_avalon_slave_read;          // mm_interconnect_0:hdmi_mm_avalon_slave_read -> hdmi_mm:s_read
	wire   [3:0] mm_interconnect_0_hdmi_mm_avalon_slave_byteenable;    // mm_interconnect_0:hdmi_mm_avalon_slave_byteenable -> hdmi_mm:s_byteenable
	wire         mm_interconnect_0_hdmi_mm_avalon_slave_readdatavalid; // hdmi_mm:s_readdatavalid -> mm_interconnect_0:hdmi_mm_avalon_slave_readdatavalid
	wire         mm_interconnect_0_hdmi_mm_avalon_slave_write;         // mm_interconnect_0:hdmi_mm_avalon_slave_write -> hdmi_mm:s_write
	wire  [31:0] mm_interconnect_0_hdmi_mm_avalon_slave_writedata;     // mm_interconnect_0:hdmi_mm_avalon_slave_writedata -> hdmi_mm:s_writedata
	wire   [0:0] mm_interconnect_0_hdmi_mm_avalon_slave_burstcount;    // mm_interconnect_0:hdmi_mm_avalon_slave_burstcount -> hdmi_mm:s_burstcount

	hdmi_mm #(
		.horz_front_porch (18),
		.horz_sync        (60),
		.horz_back_porch  (112),
		.horz_pix         (1024),
		.vert_front_porch (18),
		.vert_sync        (60),
		.vert_back_porch  (112),
		.vert_pix         (600)
	) hdmi_mm (
		.clk             (clk_clk),                                              //        clock.clk
		.reset           (~reset_reset_n),                                       //        reset.reset
		.clk_mm          (hdmi_clk_mm),                                          //      hdmi_mm.clk_mm
		.clk_pix_p       (hdmi_clk_pix_p),                                       //             .clk_pix_p
		.clk_pix_n       (hdmi_clk_pix_n),                                       //             .clk_pix_n
		.red_p           (hdmi_red_p),                                           //             .red_p
		.red_n           (hdmi_red_n),                                           //             .red_n
		.green_p         (hdmi_green_p),                                         //             .green_p
		.green_n         (hdmi_green_n),                                         //             .green_n
		.blue_p          (hdmi_blue_p),                                          //             .blue_p
		.blue_n          (hdmi_blue_n),                                          //             .blue_n
		.x               (hdmi_x),                                               //             .x
		.y               (hdmi_y),                                               //             .y
		.horz            (hdmi_horz),                                            //             .horz
		.vert            (hdmi_vert),                                            //             .vert
		.s_read          (mm_interconnect_0_hdmi_mm_avalon_slave_read),          // avalon_slave.read
		.s_write         (mm_interconnect_0_hdmi_mm_avalon_slave_write),         //             .write
		.s_address       (mm_interconnect_0_hdmi_mm_avalon_slave_address),       //             .address
		.s_writedata     (mm_interconnect_0_hdmi_mm_avalon_slave_writedata),     //             .writedata
		.s_burstcount    (mm_interconnect_0_hdmi_mm_avalon_slave_burstcount),    //             .burstcount
		.s_byteenable    (mm_interconnect_0_hdmi_mm_avalon_slave_byteenable),    //             .byteenable
		.s_waitrequest   (mm_interconnect_0_hdmi_mm_avalon_slave_waitrequest),   //             .waitrequest
		.s_readdatavalid (mm_interconnect_0_hdmi_mm_avalon_slave_readdatavalid), //             .readdatavalid
		.s_readdata      (mm_interconnect_0_hdmi_mm_avalon_slave_readdata),      //             .readdata
		.clk_x10         (clk_x10_clk)                                           //      clk_x10.clk
	);

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (32),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (4),
		.AV_BURSTCOUNT_W            (1),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (1),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (1),
		.AV_BURST_LINEWRAP          (1),
		.AV_BURST_BNDR_ONLY         (1),
		.AV_MAX_PENDING_READS       (0),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (1),
		.AV_READ_WAIT_TIME          (1),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (0)
	) master_bfm (
		.clk                    (clk_clk),                     //       clk.clk
		.reset                  (~reset_reset_n),              // clk_reset.reset
		.avm_address            (master_bfm_m0_address),       //        m0.address
		.avm_burstcount         (master_bfm_m0_burstcount),    //          .burstcount
		.avm_readdata           (master_bfm_m0_readdata),      //          .readdata
		.avm_writedata          (master_bfm_m0_writedata),     //          .writedata
		.avm_waitrequest        (master_bfm_m0_waitrequest),   //          .waitrequest
		.avm_write              (master_bfm_m0_write),         //          .write
		.avm_read               (master_bfm_m0_read),          //          .read
		.avm_byteenable         (master_bfm_m0_byteenable),    //          .byteenable
		.avm_readdatavalid      (master_bfm_m0_readdatavalid), //          .readdatavalid
		.avm_begintransfer      (),                            // (terminated)
		.avm_beginbursttransfer (),                            // (terminated)
		.avm_arbiterlock        (),                            // (terminated)
		.avm_lock               (),                            // (terminated)
		.avm_debugaccess        (),                            // (terminated)
		.avm_transactionid      (),                            // (terminated)
		.avm_readid             (8'b00000000),                 // (terminated)
		.avm_writeid            (8'b00000000),                 // (terminated)
		.avm_clken              (),                            // (terminated)
		.avm_response           (2'b00),                       // (terminated)
		.avm_writeresponsevalid (1'b0),                        // (terminated)
		.avm_readresponse       (8'b00000000),                 // (terminated)
		.avm_writeresponse      (8'b00000000)                  // (terminated)
	);

	hdmi_qsys_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                    (clk_clk),                                              //                                  clk_0_clk.clk
		.master_bfm_clk_reset_reset_bridge_in_reset_reset (~reset_reset_n),                                       // master_bfm_clk_reset_reset_bridge_in_reset.reset
		.master_bfm_m0_address                            (master_bfm_m0_address),                                //                              master_bfm_m0.address
		.master_bfm_m0_waitrequest                        (master_bfm_m0_waitrequest),                            //                                           .waitrequest
		.master_bfm_m0_burstcount                         (master_bfm_m0_burstcount),                             //                                           .burstcount
		.master_bfm_m0_byteenable                         (master_bfm_m0_byteenable),                             //                                           .byteenable
		.master_bfm_m0_read                               (master_bfm_m0_read),                                   //                                           .read
		.master_bfm_m0_readdata                           (master_bfm_m0_readdata),                               //                                           .readdata
		.master_bfm_m0_readdatavalid                      (master_bfm_m0_readdatavalid),                          //                                           .readdatavalid
		.master_bfm_m0_write                              (master_bfm_m0_write),                                  //                                           .write
		.master_bfm_m0_writedata                          (master_bfm_m0_writedata),                              //                                           .writedata
		.hdmi_mm_avalon_slave_address                     (mm_interconnect_0_hdmi_mm_avalon_slave_address),       //                       hdmi_mm_avalon_slave.address
		.hdmi_mm_avalon_slave_write                       (mm_interconnect_0_hdmi_mm_avalon_slave_write),         //                                           .write
		.hdmi_mm_avalon_slave_read                        (mm_interconnect_0_hdmi_mm_avalon_slave_read),          //                                           .read
		.hdmi_mm_avalon_slave_readdata                    (mm_interconnect_0_hdmi_mm_avalon_slave_readdata),      //                                           .readdata
		.hdmi_mm_avalon_slave_writedata                   (mm_interconnect_0_hdmi_mm_avalon_slave_writedata),     //                                           .writedata
		.hdmi_mm_avalon_slave_burstcount                  (mm_interconnect_0_hdmi_mm_avalon_slave_burstcount),    //                                           .burstcount
		.hdmi_mm_avalon_slave_byteenable                  (mm_interconnect_0_hdmi_mm_avalon_slave_byteenable),    //                                           .byteenable
		.hdmi_mm_avalon_slave_readdatavalid               (mm_interconnect_0_hdmi_mm_avalon_slave_readdatavalid), //                                           .readdatavalid
		.hdmi_mm_avalon_slave_waitrequest                 (mm_interconnect_0_hdmi_mm_avalon_slave_waitrequest)    //                                           .waitrequest
	);

endmodule
