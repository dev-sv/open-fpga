
module hdmi_qsys (
	clk_clk,
	hdmi_clk_pix_p,
	hdmi_clk_pix_n,
	hdmi_red_p,
	hdmi_red_n,
	hdmi_green_p,
	hdmi_green_n,
	hdmi_blue_p,
	hdmi_blue_n,
	memory_mem_a,
	memory_mem_ba,
	memory_mem_ck,
	memory_mem_ck_n,
	memory_mem_cke,
	memory_mem_cs_n,
	memory_mem_ras_n,
	memory_mem_cas_n,
	memory_mem_we_n,
	memory_mem_reset_n,
	memory_mem_dq,
	memory_mem_dqs,
	memory_mem_dqs_n,
	memory_mem_odt,
	memory_mem_dm,
	memory_oct_rzqin,
	pll_0_locked_export);	

	input		clk_clk;
	output		hdmi_clk_pix_p;
	output		hdmi_clk_pix_n;
	output		hdmi_red_p;
	output		hdmi_red_n;
	output		hdmi_green_p;
	output		hdmi_green_n;
	output		hdmi_blue_p;
	output		hdmi_blue_n;
	output	[14:0]	memory_mem_a;
	output	[2:0]	memory_mem_ba;
	output		memory_mem_ck;
	output		memory_mem_ck_n;
	output		memory_mem_cke;
	output		memory_mem_cs_n;
	output		memory_mem_ras_n;
	output		memory_mem_cas_n;
	output		memory_mem_we_n;
	output		memory_mem_reset_n;
	inout	[31:0]	memory_mem_dq;
	inout	[3:0]	memory_mem_dqs;
	inout	[3:0]	memory_mem_dqs_n;
	output		memory_mem_odt;
	output	[3:0]	memory_mem_dm;
	input		memory_oct_rzqin;
	output		pll_0_locked_export;
endmodule
