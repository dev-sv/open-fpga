


module tb_top(input n);


endmodule
