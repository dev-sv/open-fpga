// hdmi_qsys.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module hdmi_qsys (
		input  wire        clk_clk,        //     clk.clk
		input  wire        clk_pix_clk,    // clk_pix.clk
		input  wire        clk_x10_clk,    // clk_x10.clk
		output wire        hdmi_blue_n,    //    hdmi.blue_n
		output wire        hdmi_blue_p,    //        .blue_p
		output wire        hdmi_clk_pix_n, //        .clk_pix_n
		output wire        hdmi_clk_pix_p, //        .clk_pix_p
		output wire        hdmi_green_n,   //        .green_n
		output wire        hdmi_green_p,   //        .green_p
		output wire        hdmi_red_n,     //        .red_n
		output wire        hdmi_red_p,     //        .red_p
		output wire [10:0] hdmi_x,         //        .x
		output wire [10:0] hdmi_y,         //        .y
		output wire [10:0] hdmi_horz,      //        .horz
		output wire [10:0] hdmi_vert,      //        .vert
		output wire        hdmi_clk_st,    //        .clk_st
		input  wire        reset_reset,    //   reset.reset
		input  wire [23:0] st_in_data,     //   st_in.data
		output wire        st_in_ready,    //        .ready
		input  wire        st_in_valid     //        .valid
	);

	hdmi_st #(
		.horz_front_porch (18),
		.horz_sync        (60),
		.horz_back_porch  (112),
		.horz_pix         (1024),
		.vert_front_porch (18),
		.vert_sync        (60),
		.vert_back_porch  (112),
		.vert_pix         (600)
	) hdmi (
		.clk       (clk_clk),        //       clock.clk
		.reset     (reset_reset),    //       reset.reset
		.data      (st_in_data),     // avalon_sink.data
		.ready     (st_in_ready),    //            .ready
		.valid     (st_in_valid),    //            .valid
		.blue_n    (hdmi_blue_n),    //      hdmi_1.blue_n
		.blue_p    (hdmi_blue_p),    //            .blue_p
		.clk_pix_n (hdmi_clk_pix_n), //            .clk_pix_n
		.clk_pix_p (hdmi_clk_pix_p), //            .clk_pix_p
		.green_n   (hdmi_green_n),   //            .green_n
		.green_p   (hdmi_green_p),   //            .green_p
		.red_n     (hdmi_red_n),     //            .red_n
		.red_p     (hdmi_red_p),     //            .red_p
		.x         (hdmi_x),         //            .x
		.y         (hdmi_y),         //            .y
		.horz      (hdmi_horz),      //            .horz
		.vert      (hdmi_vert),      //            .vert
		.clk_st    (hdmi_clk_st),    //            .clk_st
		.clk_pix   (clk_pix_clk),    //     clk_pix.clk
		.clk_x10   (clk_x10_clk)     //     clk_x10.clk
	);

endmodule
