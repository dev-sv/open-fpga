// sdram_qsys.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module sdram_qsys (
		input  wire        clk_clk,       //   clk.clk
		input  wire        reset_reset_n, // reset.reset_n
		inout  wire [15:0] sdram_dq,      // sdram.dq
		output wire [11:0] sdram_address, //      .address
		output wire [1:0]  sdram_ba,      //      .ba
		output wire [1:0]  sdram_dqm,     //      .dqm
		output wire        sdram_osc,     //      .osc
		output wire        sdram_cs,      //      .cs
		output wire        sdram_we,      //      .we
		output wire        sdram_ras,     //      .ras
		output wire        sdram_cas      //      .cas
	);

	wire  [15:0] master_bfm_m0_readdata;                                 // mm_interconnect_0:master_bfm_m0_readdata -> master_bfm:avm_readdata
	wire         master_bfm_m0_waitrequest;                              // mm_interconnect_0:master_bfm_m0_waitrequest -> master_bfm:avm_waitrequest
	wire  [21:0] master_bfm_m0_address;                                  // master_bfm:avm_address -> mm_interconnect_0:master_bfm_m0_address
	wire         master_bfm_m0_read;                                     // master_bfm:avm_read -> mm_interconnect_0:master_bfm_m0_read
	wire   [1:0] master_bfm_m0_byteenable;                               // master_bfm:avm_byteenable -> mm_interconnect_0:master_bfm_m0_byteenable
	wire         master_bfm_m0_readdatavalid;                            // mm_interconnect_0:master_bfm_m0_readdatavalid -> master_bfm:avm_readdatavalid
	wire  [15:0] master_bfm_m0_writedata;                                // master_bfm:avm_writedata -> mm_interconnect_0:master_bfm_m0_writedata
	wire         master_bfm_m0_write;                                    // master_bfm:avm_write -> mm_interconnect_0:master_bfm_m0_write
	wire   [8:0] master_bfm_m0_burstcount;                               // master_bfm:avm_burstcount -> mm_interconnect_0:master_bfm_m0_burstcount
	wire  [15:0] mm_interconnect_0_sdram_avl_avalon_slave_readdata;      // sdram_avl:s_readdata -> mm_interconnect_0:sdram_avl_avalon_slave_readdata
	wire         mm_interconnect_0_sdram_avl_avalon_slave_waitrequest;   // sdram_avl:s_waitrequest -> mm_interconnect_0:sdram_avl_avalon_slave_waitrequest
	wire  [21:0] mm_interconnect_0_sdram_avl_avalon_slave_address;       // mm_interconnect_0:sdram_avl_avalon_slave_address -> sdram_avl:s_address
	wire         mm_interconnect_0_sdram_avl_avalon_slave_read;          // mm_interconnect_0:sdram_avl_avalon_slave_read -> sdram_avl:s_read
	wire   [1:0] mm_interconnect_0_sdram_avl_avalon_slave_byteenable;    // mm_interconnect_0:sdram_avl_avalon_slave_byteenable -> sdram_avl:s_byteenable
	wire         mm_interconnect_0_sdram_avl_avalon_slave_readdatavalid; // sdram_avl:s_readdatavalid -> mm_interconnect_0:sdram_avl_avalon_slave_readdatavalid
	wire         mm_interconnect_0_sdram_avl_avalon_slave_write;         // mm_interconnect_0:sdram_avl_avalon_slave_write -> sdram_avl:s_write
	wire  [15:0] mm_interconnect_0_sdram_avl_avalon_slave_writedata;     // mm_interconnect_0:sdram_avl_avalon_slave_writedata -> sdram_avl:s_writedata
	wire   [8:0] mm_interconnect_0_sdram_avl_avalon_slave_burstcount;    // mm_interconnect_0:sdram_avl_avalon_slave_burstcount -> sdram_avl:s_burstcount
	wire         rst_controller_reset_out_reset;                         // rst_controller:reset_out -> [master_bfm:reset, mm_interconnect_0:master_bfm_clk_reset_reset_bridge_in_reset_reset, sdram_avl:reset]

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (22),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (2),
		.AV_BURSTCOUNT_W            (9),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (1),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (1),
		.AV_BURST_LINEWRAP          (1),
		.AV_BURST_BNDR_ONLY         (1),
		.AV_MAX_PENDING_READS       (4),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (1),
		.AV_READ_WAIT_TIME          (1),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (0)
	) master_bfm (
		.clk                    (clk_clk),                        //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.avm_address            (master_bfm_m0_address),          //        m0.address
		.avm_burstcount         (master_bfm_m0_burstcount),       //          .burstcount
		.avm_readdata           (master_bfm_m0_readdata),         //          .readdata
		.avm_writedata          (master_bfm_m0_writedata),        //          .writedata
		.avm_waitrequest        (master_bfm_m0_waitrequest),      //          .waitrequest
		.avm_write              (master_bfm_m0_write),            //          .write
		.avm_read               (master_bfm_m0_read),             //          .read
		.avm_byteenable         (master_bfm_m0_byteenable),       //          .byteenable
		.avm_readdatavalid      (master_bfm_m0_readdatavalid),    //          .readdatavalid
		.avm_begintransfer      (),                               // (terminated)
		.avm_beginbursttransfer (),                               // (terminated)
		.avm_arbiterlock        (),                               // (terminated)
		.avm_lock               (),                               // (terminated)
		.avm_debugaccess        (),                               // (terminated)
		.avm_transactionid      (),                               // (terminated)
		.avm_readid             (8'b00000000),                    // (terminated)
		.avm_writeid            (8'b00000000),                    // (terminated)
		.avm_clken              (),                               // (terminated)
		.avm_response           (2'b00),                          // (terminated)
		.avm_writeresponsevalid (1'b0),                           // (terminated)
		.avm_readresponse       (8'b00000000),                    // (terminated)
		.avm_writeresponse      (8'b00000000)                     // (terminated)
	);

	sdram #(
		.WRITE_RECOVERY_TIME      (2),
		.PRECHARGE_COMMAND_PERIOD (2),
		.AUTO_REFRESH_PERIOD      (7),
		.LOAD_MODE_REGISTER       (3),
		.ACTIVE_READ_WRITE        (2),
		.REFRESH_PERIOD           (6400000)
	) sdram_avl (
		.clk             (clk_clk),                                                //        clock.clk
		.reset           (rst_controller_reset_out_reset),                         //        reset.reset
		.dq              (sdram_dq),                                               //        sdram.dq
		.address         (sdram_address),                                          //             .address
		.ba              (sdram_ba),                                               //             .ba
		.dqm             (sdram_dqm),                                              //             .dqm
		.osc             (sdram_osc),                                              //             .osc
		.cs              (sdram_cs),                                               //             .cs
		.we              (sdram_we),                                               //             .we
		.ras             (sdram_ras),                                              //             .ras
		.cas             (sdram_cas),                                              //             .cas
		.s_read          (mm_interconnect_0_sdram_avl_avalon_slave_read),          // avalon_slave.read
		.s_write         (mm_interconnect_0_sdram_avl_avalon_slave_write),         //             .write
		.s_address       (mm_interconnect_0_sdram_avl_avalon_slave_address),       //             .address
		.s_writedata     (mm_interconnect_0_sdram_avl_avalon_slave_writedata),     //             .writedata
		.s_burstcount    (mm_interconnect_0_sdram_avl_avalon_slave_burstcount),    //             .burstcount
		.s_byteenable    (mm_interconnect_0_sdram_avl_avalon_slave_byteenable),    //             .byteenable
		.s_waitrequest   (mm_interconnect_0_sdram_avl_avalon_slave_waitrequest),   //             .waitrequest
		.s_readdatavalid (mm_interconnect_0_sdram_avl_avalon_slave_readdatavalid), //             .readdatavalid
		.s_readdata      (mm_interconnect_0_sdram_avl_avalon_slave_readdata)       //             .readdata
	);

	sdram_qsys_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                    (clk_clk),                                                //                                  clk_0_clk.clk
		.master_bfm_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                         // master_bfm_clk_reset_reset_bridge_in_reset.reset
		.master_bfm_m0_address                            (master_bfm_m0_address),                                  //                              master_bfm_m0.address
		.master_bfm_m0_waitrequest                        (master_bfm_m0_waitrequest),                              //                                           .waitrequest
		.master_bfm_m0_burstcount                         (master_bfm_m0_burstcount),                               //                                           .burstcount
		.master_bfm_m0_byteenable                         (master_bfm_m0_byteenable),                               //                                           .byteenable
		.master_bfm_m0_read                               (master_bfm_m0_read),                                     //                                           .read
		.master_bfm_m0_readdata                           (master_bfm_m0_readdata),                                 //                                           .readdata
		.master_bfm_m0_readdatavalid                      (master_bfm_m0_readdatavalid),                            //                                           .readdatavalid
		.master_bfm_m0_write                              (master_bfm_m0_write),                                    //                                           .write
		.master_bfm_m0_writedata                          (master_bfm_m0_writedata),                                //                                           .writedata
		.sdram_avl_avalon_slave_address                   (mm_interconnect_0_sdram_avl_avalon_slave_address),       //                     sdram_avl_avalon_slave.address
		.sdram_avl_avalon_slave_write                     (mm_interconnect_0_sdram_avl_avalon_slave_write),         //                                           .write
		.sdram_avl_avalon_slave_read                      (mm_interconnect_0_sdram_avl_avalon_slave_read),          //                                           .read
		.sdram_avl_avalon_slave_readdata                  (mm_interconnect_0_sdram_avl_avalon_slave_readdata),      //                                           .readdata
		.sdram_avl_avalon_slave_writedata                 (mm_interconnect_0_sdram_avl_avalon_slave_writedata),     //                                           .writedata
		.sdram_avl_avalon_slave_burstcount                (mm_interconnect_0_sdram_avl_avalon_slave_burstcount),    //                                           .burstcount
		.sdram_avl_avalon_slave_byteenable                (mm_interconnect_0_sdram_avl_avalon_slave_byteenable),    //                                           .byteenable
		.sdram_avl_avalon_slave_readdatavalid             (mm_interconnect_0_sdram_avl_avalon_slave_readdatavalid), //                                           .readdatavalid
		.sdram_avl_avalon_slave_waitrequest               (mm_interconnect_0_sdram_avl_avalon_slave_waitrequest)    //                                           .waitrequest
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
