


module tb_top(input bit n);


endmodule
