//----------------------------------------------------------------------------------------------------
// This is the top file of the example test for Avalon Streaming BFM user guide
// The Qsys test bench system and the test program are instantiated.
//----------------------------------------------------------------------------------------------------

module top ();

	hdmi_qsys_tb tb();
    
	tb_hdmi tst();

endmodule
